.title Common Emitter Amplifier
* Model of a common emitter amplifier with a general BJT
.model QMOD	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=50 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
Q1 out bin e QMOD
C1 bin in 0.1u
R1 vcc bin 110k
R2 bin GND 10k
R4 e GND 1k
R3 vcc out 10k
VCC vcc 0 20
Vin in 0 dc 0 ac 0 SIN(0.5 0.25 1k)

.control
* tran 10u 10m
* plot v(in) v(out)
.endc

.end