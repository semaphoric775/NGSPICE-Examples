.title Pulse Generator
* First BJT Pulse Generator in AoE
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
Q1 Net-_C1-Pad2_ Net-_Q1-Pad2_ 0 Q2N3904
Q2 out Net-_C1-Pad1_ 0 Q2N3904
R1 Net-_Q1-Pad2_ in 10k
Vin in 0 dc 0 ac 0 PWL(0 0 0.0999u 0 0.1u 5)
VCC vcc 0 5
R2 vcc Net-_C1-Pad2_ 1k
R4 vcc out 1k
R3 vcc Net-_C1-Pad1_ 10k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 10n
.control
tran 10u 1m
plot v(in) v(out)
.endc

.end